`ifndef OPERATION_SVH_
`define OPERATION_SVH_

`define MMU_READ(DRIVER, ADDR, BURST, SIZE) \
	DRIVER``_ADDR <= ADDR; \
	DRIVER``_BURST <= BURST; \
	DRIVER``_SIZE <= SIZE; \
	DRIVER``_WRITE <= 1'b0; \
	DRIVER``_CLAIM <= 1'b1;

`define MMU_WRITE(DRIVER, ADDR, WRITE, SIZE, BURST) \
	DRIVER``_ADDR <= ADDR; \
	DRIVER``_WRITE_DATA <= WRITE; \
	DRIVER``_BURST <= BURST; \
	DRIVER``_SIZE <= SIZE; \
	DRIEVR``_WRITE <= 1'b1; \
	DRIVER``_CLAIM <= 1'b1;

`define MMU_RELEASE(DRIVER) \
	DRIVER``_CLAIM <= 1'b0;

`endif
