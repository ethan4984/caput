`ifndef FREELIST_SVH_
`define FREELIST_SVH_

`define FL_CLAIM_IDLE (1 << 0)
`define FL_FREE_IDLE (1 << 1)

`define FL_INIT(CONTROL) \
	CONTROL <= `FL_CLAIM_IDLE | `FL_FREE_IDLE;

`define FL_ALLOC(CONTROL, CLAIM, AVAILABLE) \
	CONTROL <= CONTROL & ~(`FL_CLAIM_IDLE) | `FL_FREE_IDLE; \
	CLAIM <= AVAILABLE

`define FL_FREE(CONTROL, FREE, INDEX) \
	CONTROL <= CONTROL & ~(`FL_FREE_IDLE) | `FL_CLAIM_IDLE; \
	FREE <= INDEX

`endif
